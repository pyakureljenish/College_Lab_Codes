module orgate(a,b,o);
input a,b;
output o;
or or1(o,a,b);
endmodule